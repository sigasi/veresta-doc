`ifndef _pixelbuffer_svh_
`define _pixelbuffer_svh_
`ifdef notdef
// TODO "Edit included file"
//      Redefine `PIXBUF_WIDTH` from '24' to '8'. Note that in the preprocessor
//      view, you can immediately see the effect on the including file: 
//      the width of the output ports gets updated as you type.
//
//      Press **Ctrl+S** to save the file and **Alt+Left** ("Back") to
//      navigate back to the including file.
`endif
`define PIXBUF_WIDTH 24
`define PIXBUF_DEPTH 8192
`endif
